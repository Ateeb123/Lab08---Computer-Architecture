module top_module
(


);





Control_Unit Control_Unit
(


);
























